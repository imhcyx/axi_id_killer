`timescale 1ns / 1ps

module sim_top #(
    parameter   ADDR_WIDTH      = 32,
    parameter   DATA_WIDTH      = 64,
    parameter   ID_WIDTH        = 4,
    parameter   MAX_R_INFLIGHT  = 8,
    parameter   MAX_W_INFLIGHT  = 8
)(
    input                       aclk,
    input                       aresetn,

    input                       s_axi_awvalid,
    output                      s_axi_awready,
    input  [ADDR_WIDTH-1:0]     s_axi_awaddr,
    input  [ID_WIDTH-1:0]       s_axi_awid,
    input  [7:0]                s_axi_awlen,
    input  [2:0]                s_axi_awsize,
    input  [1:0]                s_axi_awburst,
    input  [0:0]                s_axi_awlock,
    input  [3:0]                s_axi_awcache,
    input  [2:0]                s_axi_awprot,
    input  [3:0]                s_axi_awqos,
    input  [3:0]                s_axi_awregion,
    input                       s_axi_arvalid,
    output                      s_axi_arready,
    input  [ADDR_WIDTH-1:0]     s_axi_araddr,
    input  [ID_WIDTH-1:0]       s_axi_arid,
    input  [7:0]                s_axi_arlen,
    input  [2:0]                s_axi_arsize,
    input  [1:0]                s_axi_arburst,
    input  [0:0]                s_axi_arlock,
    input  [3:0]                s_axi_arcache,
    input  [2:0]                s_axi_arprot,
    input  [3:0]                s_axi_arqos,
    input  [3:0]                s_axi_arregion,
    input                       s_axi_wvalid,
    output                      s_axi_wready,
    input  [DATA_WIDTH-1:0]     s_axi_wdata,
    input  [DATA_WIDTH/8-1:0]   s_axi_wstrb,
    input                       s_axi_wlast,
    output                      s_axi_bvalid,
    input                       s_axi_bready,
    output [1:0]                s_axi_bresp,
    output [ID_WIDTH-1:0]       s_axi_bid,
    output                      s_axi_rvalid,
    input                       s_axi_rready,
    output [DATA_WIDTH-1:0]     s_axi_rdata,
    output [1:0]                s_axi_rresp,
    output [ID_WIDTH-1:0]       s_axi_rid,
    output                      s_axi_rlast,

    output                      m_axi_awvalid,
    input                       m_axi_awready,
    output [ADDR_WIDTH-1:0]     m_axi_awaddr,
    input                       m_axi_awid,
    output [7:0]                m_axi_awlen,
    output [2:0]                m_axi_awsize,
    output [1:0]                m_axi_awburst,
    output [0:0]                m_axi_awlock,
    output [3:0]                m_axi_awcache,
    output [2:0]                m_axi_awprot,
    output [3:0]                m_axi_awqos,
    output [3:0]                m_axi_awregion,
    output                      m_axi_arvalid,
    input                       m_axi_arready,
    output [ADDR_WIDTH-1:0]     m_axi_araddr,
    input                       m_axi_arid,
    output [7:0]                m_axi_arlen,
    output [2:0]                m_axi_arsize,
    output [1:0]                m_axi_arburst,
    output [0:0]                m_axi_arlock,
    output [3:0]                m_axi_arcache,
    output [2:0]                m_axi_arprot,
    output [3:0]                m_axi_arqos,
    output [3:0]                m_axi_arregion,
    output                      m_axi_wvalid,
    input                       m_axi_wready,
    output [DATA_WIDTH-1:0]     m_axi_wdata,
    output [DATA_WIDTH/8-1:0]   m_axi_wstrb,
    output                      m_axi_wlast,
    input                       m_axi_bvalid,
    output                      m_axi_bready,
    input  [1:0]                m_axi_bresp,
    input                       m_axi_bid,
    input                       m_axi_rvalid,
    output                      m_axi_rready,
    input  [DATA_WIDTH-1:0]     m_axi_rdata,
    input  [1:0]                m_axi_rresp,
    input                       m_axi_rid,
    input                       m_axi_rlast
);

    axi_id_killer #(
        .ADDR_WIDTH     (ADDR_WIDTH    ),
        .DATA_WIDTH     (DATA_WIDTH    ),
        .ID_WIDTH       (ID_WIDTH      ),
        .MAX_R_INFLIGHT (MAX_R_INFLIGHT),
        .MAX_W_INFLIGHT (MAX_W_INFLIGHT)
    ) uut (
        .aclk           (aclk),
        .aresetn        (aresetn),
        .s_axi_awvalid  (s_axi_awvalid),
        .s_axi_awready  (s_axi_awready),
        .s_axi_awaddr   (s_axi_awaddr),
        .s_axi_awid     (s_axi_awid),
        .s_axi_awlen    (s_axi_awlen),
        .s_axi_awsize   (s_axi_awsize),
        .s_axi_awburst  (s_axi_awburst),
        .s_axi_awlock   (s_axi_awlock),
        .s_axi_awcache  (s_axi_awcache),
        .s_axi_awprot   (s_axi_awprot),
        .s_axi_awqos    (s_axi_awqos),
        .s_axi_awregion (s_axi_awregion),
        .s_axi_arvalid  (s_axi_arvalid),
        .s_axi_arready  (s_axi_arready),
        .s_axi_araddr   (s_axi_araddr),
        .s_axi_arid     (s_axi_arid),
        .s_axi_arlen    (s_axi_arlen),
        .s_axi_arsize   (s_axi_arsize),
        .s_axi_arburst  (s_axi_arburst),
        .s_axi_arlock   (s_axi_arlock),
        .s_axi_arcache  (s_axi_arcache),
        .s_axi_arprot   (s_axi_arprot),
        .s_axi_arqos    (s_axi_arqos),
        .s_axi_arregion (s_axi_arregion),
        .s_axi_wvalid   (s_axi_wvalid),
        .s_axi_wready   (s_axi_wready),
        .s_axi_wdata    (s_axi_wdata),
        .s_axi_wstrb    (s_axi_wstrb),
        .s_axi_wlast    (s_axi_wlast),
        .s_axi_bvalid   (s_axi_bvalid),
        .s_axi_bready   (s_axi_bready),
        .s_axi_bresp    (s_axi_bresp),
        .s_axi_bid      (s_axi_bid),
        .s_axi_rvalid   (s_axi_rvalid),
        .s_axi_rready   (s_axi_rready),
        .s_axi_rdata    (s_axi_rdata),
        .s_axi_rresp    (s_axi_rresp),
        .s_axi_rid      (s_axi_rid),
        .s_axi_rlast    (s_axi_rlast),
        .m_axi_awvalid  (m_axi_awvalid),
        .m_axi_awready  (m_axi_awready),
        .m_axi_awaddr   (m_axi_awaddr),
        .m_axi_awlen    (m_axi_awlen),
        .m_axi_awsize   (m_axi_awsize),
        .m_axi_awburst  (m_axi_awburst),
        .m_axi_awlock   (m_axi_awlock),
        .m_axi_awcache  (m_axi_awcache),
        .m_axi_awprot   (m_axi_awprot),
        .m_axi_awqos    (m_axi_awqos),
        .m_axi_awregion (m_axi_awregion),
        .m_axi_arvalid  (m_axi_arvalid),
        .m_axi_arready  (m_axi_arready),
        .m_axi_araddr   (m_axi_araddr),
        .m_axi_arlen    (m_axi_arlen),
        .m_axi_arsize   (m_axi_arsize),
        .m_axi_arburst  (m_axi_arburst),
        .m_axi_arlock   (m_axi_arlock),
        .m_axi_arcache  (m_axi_arcache),
        .m_axi_arprot   (m_axi_arprot),
        .m_axi_arqos    (m_axi_arqos),
        .m_axi_arregion (m_axi_arregion),
        .m_axi_wvalid   (m_axi_wvalid),
        .m_axi_wready   (m_axi_wready),
        .m_axi_wdata    (m_axi_wdata),
        .m_axi_wstrb    (m_axi_wstrb),
        .m_axi_wlast    (m_axi_wlast),
        .m_axi_bvalid   (m_axi_bvalid),
        .m_axi_bready   (m_axi_bready),
        .m_axi_bresp    (m_axi_bresp),
        .m_axi_rvalid   (m_axi_rvalid),
        .m_axi_rready   (m_axi_rready),
        .m_axi_rdata    (m_axi_rdata),
        .m_axi_rresp    (m_axi_rresp),
        .m_axi_rlast    (m_axi_rlast)
    );

    assign m_axi_awid = 0;
    assign m_axi_arid = 0;

    initial begin
        $dumpfile("dump.vcd");
        $dumpvars;
    end

endmodule